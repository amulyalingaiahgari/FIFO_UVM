package fifo_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "transaction.sv"
  `include "driver.sv"
  `include "monitor.sv"
  `include "agent.sv"
  `include "scoreboard.sv"
  `include "environment.sv"
  `include "basic_test_seq.sv"
  `include "base_test.sv"
endpackage
